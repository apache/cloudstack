conectix             <�tap           @      @  �   ���R������G�.j���!                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������             2    ���E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                        tdbatmap      
      ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    conectix             <�tap           @      @  �   ���R������G�.j���!                                                                                                                                                                                                                                                                                                                                                                                                                                            